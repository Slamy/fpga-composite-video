`define PAL_CHROMA_B0 5
`define PAL_CHROMA_B1 0
`define PAL_CHROMA_B2 -5
`define PAL_CHROMA_A0 32
`define PAL_CHROMA_A1 -45
`define PAL_CHROMA_A2 22
`define PAL_CHROMA_B_AFTER_DOT 5
`define PAL_CHROMA_A_AFTER_DOT 5

`define NTSC_CHROMA_B0 5
`define NTSC_CHROMA_B1 0
`define NTSC_CHROMA_B2 -5
`define NTSC_CHROMA_A0 32
`define NTSC_CHROMA_A1 -48
`define NTSC_CHROMA_A2 22
`define NTSC_CHROMA_B_AFTER_DOT 5
`define NTSC_CHROMA_A_AFTER_DOT 5

`define PAL_LUMA_LOWPASS_B0 20
`define PAL_LUMA_LOWPASS_B1 41
`define PAL_LUMA_LOWPASS_B2 20
`define PAL_LUMA_LOWPASS_A0 1024
`define PAL_LUMA_LOWPASS_A1 -1530
`define PAL_LUMA_LOWPASS_A2 587
`define PAL_LUMA_LOWPASS_B_AFTER_DOT 10
`define PAL_LUMA_LOWPASS_A_AFTER_DOT 10

`define SECAM_AMPLITUDE_LOWPASS_B0 65
`define SECAM_AMPLITUDE_LOWPASS_B1 65
`define SECAM_AMPLITUDE_LOWPASS_B2 0
`define SECAM_AMPLITUDE_LOWPASS_A0 256
`define SECAM_AMPLITUDE_LOWPASS_A1 -240
`define SECAM_AMPLITUDE_LOWPASS_A2 0
`define SECAM_AMPLITUDE_LOWPASS_B_AFTER_DOT 11
`define SECAM_AMPLITUDE_LOWPASS_A_AFTER_DOT 8

`define SECAM_CHROMA_LOWPASS_B0 161
`define SECAM_CHROMA_LOWPASS_B1 161
`define SECAM_CHROMA_LOWPASS_B2 0
`define SECAM_CHROMA_LOWPASS_A0 256
`define SECAM_CHROMA_LOWPASS_A1 -216
`define SECAM_CHROMA_LOWPASS_A2 0
`define SECAM_CHROMA_LOWPASS_B_AFTER_DOT 11
`define SECAM_CHROMA_LOWPASS_A_AFTER_DOT 8

`define SECAM_PREEMPHASIS_B0 39
`define SECAM_PREEMPHASIS_B1 39
`define SECAM_PREEMPHASIS_B2 0
`define SECAM_PREEMPHASIS_A0 256
`define SECAM_PREEMPHASIS_A1 -246
`define SECAM_PREEMPHASIS_A2 0
`define SECAM_PREEMPHASIS_B_AFTER_DOT 11
`define SECAM_PREEMPHASIS_A_AFTER_DOT 8

`define CLK_PERIOD_USEC 0.020833333333333332  // .8

`define SECAM_CHROMA_DB_DDS_INCREMENT 51'd199378108503381
`define SECAM_CHROMA_DR_DDS_INCREMENT 51'd206708655146849
`define PAL_CHROMA_DDS_INCREMENT 51'd207992122400030
`define NTSC_CHROMA_DDS_INCREMENT 51'd167925390918291

`define PAL_BURST_U -8
`define PAL_BURST_V 8
`define NTSC_BURST_U -14
`define NTSC_BURST_V 4


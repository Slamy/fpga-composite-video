
`define CONFIG_SECAM_ENABLED
`define CONFIG_PAL_NTSC_ENABLED

// Optimized for YCbCr
`define CONFIG_PAL_Y_SCALER 125
`define CONFIG_PAL_U_SCALER 10
`define CONFIG_PAL_V_SCALER 15

`define CONFIG_NTSC_Y_SCALER 125
`define CONFIG_NTSC_U_SCALER 10
`define CONFIG_NTSC_V_SCALER 15

`define CONFIG_SECAM_Y_SCALER 125
`define CONFIG_SECAM_U_SCALER 10
`define CONFIG_SECAM_V_SCALER 14

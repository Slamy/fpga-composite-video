
`define CONFIG_SECAM_ENABLED
`define CONFIG_PAL_NTSC_ENABLED


`define CONFIG_SECAM_ENABLED
`define CONFIG_PAL_NTSC_ENABLED
// `define CONFIG_PAL_NTSC_CHROMA_LOWPASS

// Optimized for YCbCr
`define CONFIG_PAL_Y_SCALER 125
`define CONFIG_PAL_U_SCALER 38
`define CONFIG_PAL_V_SCALER 54

`define CONFIG_NTSC_Y_SCALER 125
`define CONFIG_NTSC_U_SCALER 38
`define CONFIG_NTSC_V_SCALER 54

`define CONFIG_SECAM_Y_SCALER 125
`define CONFIG_SECAM_U_SCALER 31
`define CONFIG_SECAM_V_SCALER 44

`define CONFIG_SECAM_DB_SWING 52
`define CONFIG_SECAM_DR_SWING 42
